netcdf pism_overrides {
    variables:
    byte pism_overrides;

    pism_overrides:air_temp_all_precip_as_snow = 272.15;
    pism_overrides:air_temp_all_precip_as_snow_doc = "Kelvin; threshold temperature below which all precipitation is snow";

    pism_overrides:air_temp_all_precip_as_rain = 274.15;
    pism_overrides:air_temp_all_precip_as_rain_doc = "Kelvin; threshold temperature above which all precipitation is rain; must exceed air_temp_all_precip_as_snow to avoid division by zero, because difference is in a denominator";

    pism_overrides:pdd_refreeze_ice_melt = "no";
    pism_overrides:pdd_refreeze_ice_melt_doc = "If set to 'yes', refreeze pdd_refreeze fraction of melted ice, otherwise all of the melted ice runs off.";

    pism_overrides:institution = "University of Alaska Fairbanks";
    pism_overrides:institution_doc = "Institution name. This string is written to output files as the 'institution' global attribute.";

    pism_overrides:backup_interval = 5.0;
    pism_overrides:backup_interval_doc = "hours; wall-clock time between automatic backups";
    
    pism_overrides:force_to_thickness_alpha = 0.05;
    pism_overrides:force_to_thickness_alpha_doc = "yr-1; exponential coefficient in force-to-thickness mechanism";

    pism_overrides:force_to_thickness_ice_free_alpha_factor = 10.0;
    pism_overrides:force_to_thickness_ice_free_alpha_factor_doc = "; force_to_thickness_alpha is multiplied by this factor in areas that are ice-free according to the target ice thickness and force_to_thickness_ice_free_thickness_threshold";


}
